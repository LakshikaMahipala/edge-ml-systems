module int8_mlp_top;
    // v0 has no I/O pins. We test int8_fc directly in TB.
endmodule
